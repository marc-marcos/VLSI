`timescale 1ns/1ps

module alu_4bit_tb;

    // TO FILL BY THE STUDENT

endmodule
